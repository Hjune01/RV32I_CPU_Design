`timescale 1ns / 1ps

module ROM (
    input  logic [31:0] addr,
    output logic [31:0] data
);
    logic [31:0] rom[0:2**8-1];

    initial begin
        //  $readmemh("code.mem", rom);

        /***************************** R-Type ***********************************/
        //rom[x]=32'b func7 _ rs2 _ rs1 _ f3_  rd _  op
        rom[0] = 32'b0000000_00001_00010_000_00100_0110011;  // ADD  x4, x2, x1     # 2 + 1 = 3
        rom[1] = 32'b0100000_00011_00001_000_00101_0110011;  // SUB  x5, x1, x3     # 1 - 3 = -2
        rom[2] = 32'b0000000_00010_00011_001_00110_0110011;  // SLL  x6, x3, x2     # 3  << 2 = 12   
        rom[3] = 32'b0000000_00001_00110_101_00111_0110011;  // SRL  x7, x6, x1     # 12 >> 1 = 6

        rom[4] = 32'b0100000_00001_00101_101_01000_0110011;  // SRA  x8,  x5, x1    # -2 >>> 1 = -1
        rom[5] = 32'b0000000_00011_00101_010_01001_0110011;  // SLT  x9,  x5, x3    # (-2 < 3) ? 1 : 0 = 1
        rom[6] = 32'b0000000_00110_00111_011_01010_0110011;  // SLTU x10, x7, x6    # (6 < 12) ? 1 : 0 = 1
        rom[7] = 32'b0000000_00111_00011_100_01011_0110011;  // XOR  x11, x3, x7    # 3 ^ 6 = 5 
        rom[8] = 32'b0000000_00011_00111_110_01100_0110011;  // OR   x12, x7, x3    # 6 | 3 = 7  
        rom[9] = 32'b0000000_01100_00110_111_01101_0110011;  // AND  x13, x6, x12   # 12 & 7 = 4
        /***************************** I-Type ***********************************/
        //rom[x]= 32'b   imm12   _ rs1 _f3 _ rd  _  op 
        rom[10] = 32'b00000001010_00111_000_01110_0010011;   // ADDI  x14, x7, 10   # 6 + 10 = 16   
        rom[11] = 32'b00000000010_00100_010_01111_0010011;   // SLTI  x15, x4, 2    # (4 < 2) ? 1 : 0 = 0
        rom[12] = 32'b00000001010_00111_011_10000_0010011;   // SLTIU x16, x7, 10   # (6 < 10) ? 1 : 0 = 1 
        rom[13] = 32'b00000000111_00110_100_10001_0010011;   // XORI  x17, x6, 7    # 12 ^ 7 = 11
        rom[14] = 32'b00000000110_10001_110_10010_0010011;   // ORI   x18, x17, 6   # 11 | 6 = 15   
        rom[15] = 32'b00000000110_10001_111_10011_0010011;   // ANDI  x19, x17, 6   # 11 & 6 = 2  
        //rom[x]= 32'b   imm12   _ rs1 _f3 _ rd  _  op          I-Type shamt
        rom[16] = 32'b00000000010_10001_001_10100_0010011;   // SLLI  x20, x17, 2   # 11 << 2 = 44
        rom[17] = 32'b00000000010_10001_101_10101_0010011;   // SRLI  x21, x17, 2   # 11 >> 2 = 2
        rom[18] = 32'b01000000010_10001_101_10110_0010011;   // SRAI  x22, x5, 1    # -2 >>> 1 = -1
        /***************************** S-Type ***********************************/
        //rom[x]=32'b  imm7  _ rs2 _ rs1 _f3 _ imm5_  op 
        rom[19] = 32'b0000000_10010_00000_010_01000_0100011;  // SW x18,  8(x0)     # 00000000_00000000_00000000_00001111 (15 저장)
        rom[20] = 32'b0000000_00101_00000_000_01010_0100011;  // SB x5,   10(x0)    # xxxxxxxx_11111110_xxxxxxxx_xxxxxxxx (-2 저장)
        rom[21] = 32'b0000000_01110_00000_001_01000_0100011;  // SH x14,  8(x0)     # xxxxxxxx_xxxxxxxx_00000000_00010000 (16 저장)
        /***************************** L-Type ***********************************/
        //rom[x]=32'b imm12      _ rs1 _f3 _ rd  _ op  
        rom[22] = 32'b000000001010_00000_000_10111_0000011;  // LB  x23, 10(x0)     # 24'b1_11111110   (-2)
        rom[23] = 32'b000000001000_00000_001_10111_0000011;  // LH  x23, 8(x0)      # 16'b0_00000000_00010000 (16)
        rom[24] = 32'b000000001000_00000_010_10111_0000011;  // LW  x23, 8(x0)      # 00000000_11111110_00000000_00010000 (16,646,160)
        rom[25] = 32'b000000001010_00000_100_10111_0000011;  // LBU x23, 10(x0)     # 24'b0_11111110   (254)
        rom[26] = 32'b000000001000_00000_101_10111_0000011;  // LHU x23, 8(x0)      # 16'b0_00000000_00010000 (16)
        /***************************** B-Type ***********************************/
        //rom[x]= 32'b imm7  _ rs2 _ rs1 _f3 _ imm5_  op         B-Type
        rom[27] = 32'b0000000_00010_00010_000_01000_1100011;  // BEQ   x2, x2, 8    # 2  = 2 
        rom[29] = 32'b0000000_00001_00010_001_01000_1100011;  // BNE   x2, x1, 8    # 2  != 1
        rom[31] = 32'b0000000_00100_00101_100_01000_1100011;  // BLT   x5, x8, 8    # -2 < -1   
        rom[33] = 32'b0000000_00101_00100_101_01000_1100011;  // BGE   x8, x5, 8    # -1 >= -2
        rom[35] = 32'b0000000_00010_00001_110_01000_1100011;  // BLTU  x1, x2, 8    # 1 < 2
        rom[37] = 32'b0000000_00001_00010_101_01000_1100011;  // BGEU  x2, x1, 8    # 2 >= 1
        /***************************** LU-Type ***********************************/
        //rom[x]= 32'b         imm20         _ rd  _   op
        rom[39] = 32'b00000_00000_00000_00101_11000_0110111;  // LUI x24, 5         # mem[24] : 5 << 12 = 20480
        /***************************** AU-Type ***********************************/
        //rom[x]= 32'b         imm20         _ rd  _   op
        rom[40] = 32'b00000_00000_00000_00101_11001_0010111;  // AUIPC x25, 5       # mem[25] : PCOutData + (5 << 12)
        /***************************** J-Type ***********************************/
        //rom[x]=32'b          imm           _ rd  _  op         J Type
        rom[41] = 32'b0_0000000100_0_00000000_11010_1101111;  // JAL x26, 8         # PC=164, mem[26] : 164 + 4 = 168, PC = 164 + 8 = 172 
        /***************************** JL-Type **********************************/
        //rom[x]= 32'b   imm12    _ rs1 _f3 _ rd  _ op           JL Type
        rom[43] = 32'b000001111000_10100_000_11011_1100111;  // JALR x27, x20, 120  # PC=172, mem[27] : 172 + 4 = 176, PC = 44(rs1) + 120(imm) = 164 

    end

    assign data = rom[addr[31:2]];
endmodule
